CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 300 9
64 124 2496 1346
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
64 124 2496 1346
144179218 256
0
6 Title:
5 Name:
0
0
0
9
11 Multimeter~
205 443 238 0 21 21
0 3 8 9 4 0 0 0 0 0
32 54 48 46 48 48 32 86 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -19 28 -11
3 MM3
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
7 Ground~
168 380 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
11 Multimeter~
205 488 178 0 21 21
0 5 10 11 3 0 0 0 0 0
32 49 48 46 48 48 48 32 0 0
0 86
0
0 0 16464 270
6 1.000u
-21 -19 21 -11
3 MM2
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
11 Multimeter~
205 512 115 0 21 21
0 5 12 13 6 0 0 0 0 0
32 50 48 46 48 48 32 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
11 Multimeter~
205 435 115 0 21 21
0 7 14 15 5 0 0 0 0 0
32 51 48 46 48 48 32 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
9 V Source~
197 401 200 0 2 5
0 7 2
0
0 0 17264 0
4 110V
10 0 38 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
7734 0 0
0
0
9 Resistor~
219 471 245 0 2 5
0 4 3
0
0 0 880 90
1 6
11 0 18 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 471 300 0 3 5
0 2 4 -1
0
0 0 880 90
1 5
11 0 18 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 541 200 0 3 5
0 2 6 -1
0
0 0 880 90
3 5.5
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
11
1 0 3 0 0 4096 0 1 0 0 7 2
459 220
471 220
4 0 4 0 0 4096 0 1 0 0 6 2
459 270
471 270
1 2 2 0 0 8192 0 2 6 0 0 3
380 219
380 221
401 221
0 2 2 0 0 8192 0 0 6 5 0 3
471 335
401 335
401 221
1 1 2 0 0 4224 0 9 8 0 0 4
541 218
541 335
471 335
471 318
1 2 4 0 0 4224 0 7 8 0 0 2
471 263
471 282
4 2 3 0 0 8320 0 3 7 0 0 3
472 210
471 210
471 227
1 0 5 0 0 4096 0 3 0 0 11 2
472 160
472 140
4 2 6 0 0 12416 0 4 9 0 0 4
537 138
537 140
541 140
541 182
1 1 7 0 0 4224 0 6 5 0 0 3
401 179
401 138
410 138
4 1 5 0 0 8320 0 5 4 0 0 4
460 138
460 140
487 140
487 138
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
9181286 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 50 2000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
