CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 0 30 300 9
0 71 2560 1078
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 2560 1078
144179218 0
0
6 Title:
5 Name:
0
0
0
16
7 Ground~
168 530 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Multimeter~
205 590 65 0 21 21
0 3 12 13 4 0 0 0 0 0
32 52 46 48 49 52 32 65 0 0
2 86
0
0 0 16464 0
7 100.00p
-24 -19 25 -11
3 MM5
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 210 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
11 Multimeter~
205 580 170 0 21 21
0 6 14 15 5 0 0 0 0 0
32 51 54 46 52 57 32 86 0 0
2 82
0
0 0 16464 782
8 100.0Meg
-28 -37 28 -29
3 MM4
-11 -47 10 -39
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
6153 0 0
0
0
11 Multimeter~
205 640 120 0 21 21
0 4 16 17 6 0 0 0 0 0
32 54 46 48 56 49 32 65 0 0
2 86
0
0 0 16464 270
6 1.000u
-21 -36 21 -28
3 MM3
-11 -46 10 -38
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
11 Multimeter~
205 680 65 0 21 21
0 4 18 19 7 0 0 0 0 0
32 56 46 48 55 56 32 65 0 0
2 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
11 Signal Gen~
195 517 155 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1134267597
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 1723754235
20
1 60 0 311.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -311/311V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 311.1 60 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
9 Inductor~
219 622 220 0 2 5
0 2 5
0
0 0 8400 90
4 0.1H
4 -4 32 4
2 L2
11 -14 25 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
10 Capacitor~
219 732 170 0 2 5
0 2 8
0
0 0 8400 90
5 100uF
5 0 40 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
10 Capacitor~
219 410 170 0 2 5
0 2 9
0
0 0 8400 90
5 100uF
4 0 39 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
9 Inductor~
219 300 170 0 2 5
0 2 10
0
0 0 8400 90
4 0.1H
4 -4 32 4
2 L1
11 -14 25 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
11 Signal Gen~
195 195 155 0 19 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1134270874
20
1 60 0 311.2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -311/311V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 311.2 60 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 622 180 0 2 5
0 5 6
0
0 0 8432 90
1 6
11 0 18 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 732 120 0 2 5
0 8 7
0
0 0 8432 90
1 5
11 0 18 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 410 120 0 2 5
0 9 11
0
0 0 8432 90
1 5
11 0 18 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 300 120 0 2 5
0 10 11
0
0 0 8432 90
1 6
11 0 18 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
19
1 1 3 0 0 4224 0 7 2 0 0 3
548 150
548 88
565 88
4 0 4 0 0 4096 0 2 0 0 7 2
615 88
624 88
1 0 2 0 0 4096 0 1 0 0 11 2
530 219
547 219
1 0 2 0 0 0 0 3 0 0 15 2
210 184
225 184
4 2 5 0 0 4224 0 4 8 0 0 2
596 202
622 202
1 4 6 0 0 4224 0 4 5 0 0 2
596 152
624 152
1 1 4 0 0 4224 0 6 5 0 0 3
655 88
624 88
624 102
2 4 6 0 0 0 0 13 5 0 0 3
622 162
624 162
624 152
4 2 7 0 0 8320 0 6 14 0 0 4
705 88
705 86
732 86
732 102
1 1 2 0 0 8336 0 9 8 0 0 4
732 179
732 250
622 250
622 238
2 1 2 0 0 0 0 7 8 0 0 5
548 160
547 160
547 250
622 250
622 238
2 1 8 0 0 4224 0 9 14 0 0 2
732 161
732 138
2 1 5 0 0 0 0 8 13 0 0 4
622 202
622 187
622 187
622 198
1 1 2 0 0 128 0 10 11 0 0 4
410 179
410 205
300 205
300 188
2 1 2 0 0 0 0 12 11 0 0 5
226 160
225 160
225 205
300 205
300 188
2 1 9 0 0 4224 0 10 15 0 0 2
410 161
410 138
2 1 10 0 0 4224 0 11 16 0 0 2
300 152
300 138
2 2 11 0 0 8320 0 15 16 0 0 4
410 102
410 86
300 86
300 102
1 2 11 0 0 0 0 12 16 0 0 5
226 150
225 150
225 86
300 86
300 102
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0833333 0.000333333 0.000333333
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
11799118 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 5000
1
517 155
0 0 0 0 0	7 0 0 0
3213960 8419392 100 100 0 0
77 66 2507 486
0 831 2560 1399
2507 66
77 66
2507 66
2507 486
0 0
0.08333 0 800 -400 0.08333 0.08333
12401 0
4 0.02 2000
1
548 111
0 3 0 0 1	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
