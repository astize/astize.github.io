CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 300 9
0 71 2560 1400
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 2560 1400
144179218 256
0
6 Title:
5 Name:
0
0
0
15
11 Multimeter~
205 433 94 0 21 21
0 3 12 13 4 0 0 0 0 0
32 55 49 52 46 51 109 65 0 0
0 86
0
0 0 16464 782
6 1.000u
-21 -19 21 -11
3 MM8
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
11 Multimeter~
205 419 40 0 21 21
0 6 14 15 3 0 0 0 0 0
45 50 46 56 53 55 32 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM7
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
11 Multimeter~
205 486 40 0 21 21
0 5 16 17 3 0 0 0 0 0
32 51 46 53 55 49 32 65 0 0
0 86
0
0 0 16464 512
6 1.000u
-21 -19 21 -11
3 MM6
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
9 V Source~
197 254 191 0 2 5
0 8 2
0
0 0 16752 512
3 20V
13 0 34 8
2 E4
17 -10 31 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
6153 0 0
0
0
9 V Source~
197 134 191 0 2 5
0 9 2
0
0 0 16752 0
3 10V
13 0 34 8
2 E3
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
5394 0 0
0
0
7 Ground~
168 115 227 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 374 226 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
9 V Source~
197 393 190 0 2 5
0 11 2
0
0 0 16752 0
3 10V
13 0 34 8
2 E1
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3747 0 0
0
0
9 V Source~
197 513 190 0 2 5
0 10 2
0
0 0 16752 512
3 20V
13 0 34 8
2 E2
17 -10 31 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3549 0 0
0
0
9 Resistor~
219 254 116 0 2 5
0 8 7
0
0 0 8432 90
1 2
11 0 18 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 134 116 0 2 5
0 9 7
0
0 0 8432 90
1 1
11 0 18 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 194 151 0 3 5
0 2 7 -1
0
0 0 8432 90
2 18
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 453 150 0 3 5
0 2 4 -1
0
0 0 8432 90
2 18
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 393 115 0 2 5
0 11 6
0
0 0 8432 90
1 1
11 0 18 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 513 115 0 2 5
0 10 5
0
0 0 8432 90
1 2
11 0 18 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
17
0 1 3 0 0 4096 0 0 1 4 0 3
452 63
452 76
449 76
2 4 4 0 0 4224 0 13 1 0 0 3
453 132
453 126
449 126
1 2 5 0 0 8320 0 3 15 0 0 3
511 63
513 63
513 97
4 4 3 0 0 4224 0 2 3 0 0 2
444 63
461 63
2 1 6 0 0 8320 0 14 2 0 0 3
393 97
394 97
394 63
0 2 7 0 0 4096 0 0 10 11 0 3
194 68
254 68
254 98
1 0 2 0 0 4096 0 6 0 0 10 2
115 221
134 221
2 0 2 0 0 8192 0 4 0 0 10 3
254 212
254 237
193 237
1 1 8 0 0 4224 0 10 4 0 0 2
254 134
254 170
2 1 2 0 0 12416 0 5 12 0 0 4
134 212
134 237
194 237
194 169
2 2 7 0 0 4224 0 12 11 0 0 5
194 133
194 68
137 68
137 98
134 98
1 1 9 0 0 4224 0 5 11 0 0 2
134 170
134 134
1 0 2 0 0 0 0 7 0 0 16 2
374 220
393 220
2 0 2 0 0 0 0 9 0 0 16 3
513 211
513 236
452 236
1 1 10 0 0 4224 0 15 9 0 0 2
513 133
513 169
2 1 2 0 0 128 0 8 13 0 0 4
393 211
393 236
453 236
453 168
1 1 11 0 0 4224 0 8 14 0 0 2
393 169
393 133
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
198922 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5 30
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
