CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 30 300 9
0 71 2560 735
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 2560 735
144179218 0
0
6 Title:
5 Name:
0
0
0
9
11 Signal Gen~
195 282 158 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1124951654
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -438896261
20
1 50 0 141.4 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -141/141V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 141.4 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
9 Inductor~
219 392 133 0 2 5
0 3 4
0
0 0 8400 270
6 31.8mH
-4 -4 38 4
2 L1
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
7 Ground~
168 316 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 520 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
11 Multimeter~
205 555 85 0 21 21
0 6 8 9 5 0 0 0 0 0
32 56 46 50 55 57 32 65 0 0
2 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
9 Inductor~
219 596 133 0 2 5
0 5 7
0
0 0 8400 270
6 31.8mH
-4 -4 38 4
2 L2
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
11 Signal Gen~
195 486 158 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1124951654
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -438896261
20
1 50 0 141.4 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -141/141V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 141.4 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
9 Resistor~
219 392 193 0 3 5
0 2 4 -1
0
0 0 8432 90
1 7
11 0 18 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 596 193 0 3 5
0 2 7 -1
0
0 0 8432 90
1 7
11 0 18 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9
1 0 2 0 0 4112 0 3 0 0 3 2
316 224
316 211
1 1 3 0 0 8336 0 1 2 0 0 4
313 153
313 108
392 108
392 115
2 1 2 0 0 8336 0 1 8 0 0 3
313 163
313 211
392 211
2 2 4 0 0 4240 0 8 2 0 0 2
392 175
392 151
1 0 2 0 0 0 0 4 0 0 8 2
520 224
520 211
4 1 5 0 0 4224 0 5 6 0 0 3
580 108
596 108
596 115
1 1 6 0 0 4224 0 7 5 0 0 3
517 153
517 108
530 108
2 1 2 0 0 128 0 7 9 0 0 3
517 163
517 211
596 211
2 2 7 0 0 4224 0 9 6 0 0 2
596 175
596 151
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
853168 1210432 100 100 0 0
0 0 0 0
113 203 274 273
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 0.1
1
517 115
0 6 0 0 1	0 7 0 0
1245668 8550464 100 100 0 0
77 66 2507 576
0 734 2560 1399
2507 66
77 66
2507 66
2507 576
0 0
0.1 0 150 -150 0.1 0.1
12401 0
4 0.03 1000
1
517 118
0 6 0 0 1	0 7 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
