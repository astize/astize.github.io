CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 300 9
0 71 2560 1400
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 2560 1400
144179218 256
0
6 Title:
5 Name:
0
0
0
25
7 Ground~
168 745 136 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 550 144 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 549 284 0 1 3
0 2
0
0 0 53360 782
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 733 173 0 1 3
0 2
0
0 0 53360 270
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 583 49 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 380 301 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 650 300 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
11 Multimeter~
205 758 224 0 21 21
0 5 14 15 2 0 0 0 0 0
32 49 46 53 48 48 32 86 0 0
0 82
0
0 0 16464 602
8 100.0Meg
-28 -19 28 -11
4 MM11
-14 -29 14 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3747 0 0
0
0
11 Multimeter~
205 721 224 0 21 21
0 5 16 17 6 0 0 0 0 0
32 53 48 46 48 48 109 65 0 0
0 86
0
0 0 16464 602
6 1.000u
-21 -19 21 -11
4 MM10
-14 -29 14 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
11 Multimeter~
205 635 58 0 21 21
0 3 18 19 7 0 0 0 0 0
32 53 48 46 48 48 109 65 0 0
0 86
0
0 0 16464 512
6 1.000u
-21 -19 21 -11
3 MM9
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
7931 0 0
0
0
11 Multimeter~
205 635 21 0 21 21
0 3 20 21 2 0 0 0 0 0
32 49 46 53 48 48 32 86 0 0
0 82
0
0 0 16464 512
8 100.0Meg
-28 -19 28 -11
3 MM8
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
9325 0 0
0
0
11 Multimeter~
205 560 223 0 21 21
0 4 22 23 8 0 0 0 0 0
32 53 48 46 48 48 109 65 0 0
0 86
0
0 0 16464 782
6 1.000u
-21 -19 21 -11
3 MM7
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
11 Multimeter~
205 524 223 0 21 21
0 4 24 25 2 0 0 0 0 0
32 49 46 53 48 48 32 86 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -19 28 -11
3 MM6
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3834 0 0
0
0
9 V Source~
197 575 155 0 2 5
0 4 2
0
0 0 16880 180
4 1.5V
14 -5 42 3
3 Vs6
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3363 0 0
0
0
9 V Source~
197 705 110 0 2 5
0 3 2
0
0 0 16752 0
4 1.5V
10 0 38 8
3 Vs5
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
7668 0 0
0
0
9 V Source~
197 665 270 0 2 5
0 5 2
0
0 0 16752 270
4 1.5V
-14 -20 14 -12
3 Vs4
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4718 0 0
0
0
9 V Source~
197 395 270 0 2 5
0 11 2
0
0 0 16752 270
4 1.5V
-14 -20 14 -12
3 Vs3
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3874 0 0
0
0
9 V Source~
197 435 110 0 2 5
0 13 9
0
0 0 16752 0
4 1.5V
10 0 38 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6671 0 0
0
0
9 V Source~
197 305 155 0 2 5
0 10 12
0
0 0 16880 0
4 1.5V
10 0 38 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3789 0 0
0
0
9 Resistor~
219 575 110 0 3 5
0 2 7 -1
0
0 0 8432 90
2 30
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 705 155 0 4 5
0 6 2 0 -1
0
0 0 8432 90
2 30
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 615 270 0 4 5
0 8 2 0 -1
0
0 0 8432 0
2 30
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 345 270 0 4 5
0 12 2 0 -1
0
0 0 8432 0
2 30
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 435 155 0 2 5
0 11 9
0
0 0 8432 90
2 30
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 305 110 0 2 5
0 10 13
0
0 0 8432 90
2 30
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
25
2 1 2 0 0 8320 0 15 1 0 0 3
705 131
705 130
745 130
2 1 2 0 0 0 0 14 2 0 0 3
575 132
550 132
550 138
1 4 2 0 0 128 0 4 8 0 0 3
740 174
741 174
741 205
1 4 2 0 0 0 0 3 13 0 0 3
542 285
540 285
540 255
1 2 2 0 0 0 0 7 16 0 0 3
650 294
650 271
643 271
1 0 3 0 0 4224 0 11 0 0 12 3
660 44
705 44
705 81
4 1 2 0 0 128 0 11 5 0 0 3
610 44
610 43
583 43
1 0 4 0 0 8320 0 13 0 0 15 3
540 205
540 185
575 185
0 1 5 0 0 4224 0 0 8 11 0 3
704 271
741 271
741 255
4 1 6 0 0 8320 0 9 21 0 0 3
704 205
705 205
705 173
1 1 5 0 0 0 0 16 9 0 0 3
685 271
704 271
704 255
1 1 3 0 0 0 0 10 15 0 0 3
660 81
705 81
705 89
4 2 7 0 0 4224 0 10 20 0 0 3
610 81
575 81
575 92
4 1 8 0 0 8320 0 12 22 0 0 3
576 255
576 270
597 270
1 1 4 0 0 0 0 12 14 0 0 3
576 205
575 205
575 174
1 2 2 0 0 128 0 6 17 0 0 4
380 295
380 285
373 285
373 271
2 1 2 0 0 128 0 14 20 0 0 2
575 132
575 128
2 2 2 0 0 128 0 15 21 0 0 2
705 131
705 137
2 2 2 0 0 128 0 22 16 0 0 3
633 270
633 271
643 271
2 2 9 0 0 4224 0 18 24 0 0 2
435 131
435 137
1 1 10 0 0 4224 0 19 25 0 0 2
305 134
305 128
1 1 11 0 0 8320 0 17 24 0 0 3
415 271
435 271
435 173
2 2 2 0 0 128 0 23 17 0 0 3
363 270
363 271
373 271
2 1 12 0 0 4224 0 19 23 0 0 3
305 176
305 270
327 270
2 1 13 0 0 8320 0 25 18 0 0 4
305 92
305 50
435 50
435 89
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2099592 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.5 1
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
