CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 300 9
0 71 2560 1400
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 2560 1400
144179218 256
0
6 Title:
5 Name:
0
0
0
10
7 Ground~
168 374 226 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Multimeter~
205 570 184 0 21 21
0 5 9 10 2 0 0 0 0 0
32 49 52 46 48 48 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -37 28 -29
3 MM4
-11 -47 10 -39
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
4441 0 0
0
0
11 Multimeter~
205 568 109 0 21 21
0 5 11 12 3 0 0 0 0 0
32 56 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 602
8 100.0Meg
-28 -37 28 -29
3 MM2
-11 -47 10 -39
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3618 0 0
0
0
11 Multimeter~
205 479 144 0 21 21
0 3 13 14 2 0 0 0 0 0
32 54 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -37 28 -29
3 MM1
-11 -47 10 -39
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
6153 0 0
0
0
11 Multimeter~
205 365 110 0 21 21
0 4 15 16 3 0 0 0 0 0
32 52 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 90
8 100.0Meg
-28 -37 28 -29
3 MM0
-11 -47 10 -39
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
5394 0 0
0
0
9 V Source~
197 393 190 0 2 5
0 4 2
0
0 0 17264 0
3 10V
13 0 34 8
2 E1
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
7734 0 0
0
0
9 V Source~
197 513 190 0 2 5
0 5 2
0
0 0 17264 512
3 14V
13 0 34 8
2 E2
17 -10 31 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
9914 0 0
0
0
9 Resistor~
219 453 150 0 3 5
0 2 3 -1
0
0 0 240 90
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 393 115 0 2 5
0 4 3
0
0 0 112 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 513 115 0 2 5
0 5 3
0
0 0 112 90
2 4k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
15
4 0 2 0 0 4096 0 4 0 0 12 2
463 176
453 176
1 0 3 0 0 4096 0 4 0 0 13 2
463 126
453 126
1 0 4 0 0 4096 0 5 0 0 14 2
382 141
393 141
4 0 3 0 0 4096 0 5 0 0 15 2
382 91
393 91
1 0 5 0 0 4096 0 3 0 0 11 2
551 140
513 140
4 0 3 0 0 4096 0 3 0 0 15 2
551 90
513 90
1 0 2 0 0 4096 0 1 0 0 12 2
374 220
393 220
1 1 5 0 0 8320 0 2 7 0 0 3
554 166
554 169
513 169
4 0 2 0 0 4096 0 2 0 0 10 2
554 216
513 216
2 0 2 0 0 8192 0 7 0 0 12 3
513 211
513 236
452 236
1 1 5 0 0 0 0 10 7 0 0 2
513 133
513 169
2 1 2 0 0 12416 0 6 8 0 0 4
393 211
393 236
453 236
453 168
2 0 3 0 0 4096 0 8 0 0 15 2
453 132
453 80
1 1 4 0 0 4224 0 6 9 0 0 2
393 169
393 133
2 2 3 0 0 8320 0 9 10 0 0 4
393 97
393 80
513 80
513 97
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3738122 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 3 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
